/*
* -----------------------------------------------------------------
* COMPANY : Ruhr University Bochum
* AUTHOR  : Amir Moradi (amir.moradi@rub.de) Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de)
* DOCUMENT: https://eprint.iacr.org/2020/
* -----------------------------------------------------------------
*
* Copyright (c) 2020, Amir Moradi, Aein Rezaei Shahmirzadi
*
* All rights reserved.
*
* THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
* ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
* WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
* DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
* DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
* (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
* LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
* ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
* (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
* SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*
* Please see LICENSE and README for license and further instructions.
*/

module GF256_INV ( clk, dcba1, dcba2, hgfe1, hgfe2, FreshRadnom, dcba1_out, 
        dcba2_out, hgfe1_out, hgfe2_out );
  (* SILVER="[3:0]_0" *)input [3:0] dcba1;
  (* SILVER="[3:0]_1" *)input [3:0] dcba2;
  (* SILVER="[7:4]_0" *) input [3:0] hgfe1;
  (* SILVER="[7:4]_1" *) input [3:0] hgfe2;
  (* SILVER="[3:0]_0" *) output [3:0] dcba1_out;
  (* SILVER="[3:0]_1" *) output [3:0] dcba2_out;
  (* SILVER="[7:4]_0" *) output [3:0] hgfe1_out;
  (* SILVER="[7:4]_1" *) output [3:0] hgfe2_out;
  (* SILVER="clock" *) input clk;
  (* SILVER="refresh" *) input FreshRadnom;
  wire   Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n47,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n46,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n45,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n44,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n43,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n42,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n41,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n40,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n39,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n38,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n37,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n36,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n35,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n34,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n33,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n32,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n31,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n30,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n29,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n28,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n27,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n26,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n25,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n24,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n23,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n22,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n21,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n20,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n19,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n18,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n17,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n16,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n15,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n14,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n13,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n12,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n11,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n10,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n9,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n8,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n7,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n6,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n5,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n4,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n3,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n2,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n1,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n46,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n45,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n44,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n43,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n42,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n41,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n40,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n39,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n38,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n37,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n36,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n35,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n34,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n33,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n32,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n31,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n30,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n29,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n28,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n27,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n26,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n25,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n24,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n23,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n22,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n21,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n20,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n19,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n18,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n17,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n16,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n15,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n11,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n10,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n9,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n8,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n7,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n6,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n5,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n4,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n3,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n2,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n1,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n49,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n48,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n47,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n46,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n45,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n44,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n43,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n42,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n41,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n40,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n39,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n38,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n37,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n36,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n35,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n34,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n33,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n32,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n31,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n30,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n29,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n28,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n27,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n26,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n17,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n16,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n15,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n14,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n13,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n12,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n11,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n10,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n9,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n8,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n7,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n6,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n5,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n4,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n3,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n2,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n1,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n44,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n43,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n42,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n41,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n40,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n39,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n38,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n37,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n36,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n35,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n34,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n33,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n32,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n31,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n30,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n29,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n28,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n27,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n26,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n25,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n24,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n23,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n22,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n21,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n20,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n19,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n18,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n17,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n16,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n15,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n14,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n13,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n12,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n11,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n10,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n9,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n8,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n7,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n6,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n5,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n4,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n3,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n2,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n1,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n12,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n11,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n10,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n9,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n8,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n7,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n6,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n5,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n4,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n3,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n2,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n1,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n34,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n33,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n32,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n31,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n30,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n29,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n28,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n27,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n26,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n25,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n24,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n23,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n22,
         Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n21,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_n3,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_n2,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_n1,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_n3,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_n2,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_n1,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n9,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n8,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n7,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n4,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n3,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n2,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n1,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n21,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n20,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n19,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n18,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n17,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n16,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n15,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n14,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n13,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n12,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n11,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n10,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n9,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n8,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n7,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n4,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n3,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n2,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n1,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n4,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n3,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n2,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n1,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n14,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n13,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n12,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n11,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n10,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n9,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n8,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n7,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n4,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n3,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n2,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n1,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n9,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n8,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n7,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n4,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n3,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n2,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n1,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n11,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n10,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n9,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n8,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n7,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n4,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n3,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n2,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n1,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n4,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n3,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n2,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n1,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n12,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n11,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n10,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n9,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n8,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n7,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n4,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n3,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n2,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n1,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n10,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n9,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n8,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n7,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n4,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n3,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n2,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n1,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n5,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n6,
         Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n5,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n90,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n89,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n143,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n142,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n141,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n140,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n152,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n151,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n150,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n149,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n148,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n147,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n146,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n145,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n144,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n143,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n142,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n141,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n140,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n140,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100,
         Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n90,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n89,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n143,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n142,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n141,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n140,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n152,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n151,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n150,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n149,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n148,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n147,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n146,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n145,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n144,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n143,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n142,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n141,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n140,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n140,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100,
         Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99;
  wire   [3:0] dcba1_reg1;
  wire   [3:0] dcba2_reg1;
  wire   [4:1] sq_scl_mul_out1;
  wire   [4:1] sq_scl_mul_out2;
  wire   [3:0] hgfe1_reg1;
  wire   [3:0] hgfe2_reg1;
  wire   [3:0] dcba1_reg2;
  wire   [3:0] dcba2_reg2;
  wire   [4:1] sq_scl_mul_out1_reg;
  wire   [4:1] sq_scl_mul_out2_reg;
  wire   [3:0] hgfe1_reg2;
  wire   [3:0] hgfe2_reg2;
  wire   [3:0] dcba1_reg3;
  wire   [3:0] dcba2_reg3;
  wire   [3:0] GF16_inv_out1;
  wire   [3:0] GF16_inv_out2;
  wire   [3:0] hgfe1_reg3;
  wire   [3:0] hgfe2_reg3;
  wire   [3:0] dcba1_reg4;
  wire   [3:0] dcba2_reg4;
  wire   [3:0] GF16_inv_out1_reg;
  wire   [3:0] GF16_inv_out2_reg;
  wire   [3:0] hgfe1_reg4;
  wire   [3:0] hgfe2_reg4;
  wire   [4:1] Inst_Gf6_sq_scl_mul_Canright_t_reg;
  wire   [4:1] Inst_Gf6_sq_scl_mul_Canright_z_reg;
  wire   [4:1] Inst_Gf6_sq_scl_mul_Canright_y_reg;
  wire   [4:1] Inst_Gf6_sq_scl_mul_Canright_x_reg;
  wire   [4:1] Inst_Gf6_sq_scl_mul_Canright_t;
  wire   [4:1] Inst_Gf6_sq_scl_mul_Canright_z;
  wire   [4:1] Inst_Gf6_sq_scl_mul_Canright_y;
  wire   [4:1] Inst_Gf6_sq_scl_mul_Canright_x;
  wire   [8:1] Inst_GF16_inv_282_t_reg;
  wire   [8:1] Inst_GF16_inv_282_z_reg;
  wire   [8:1] Inst_GF16_inv_282_y_reg;
  wire   [8:1] Inst_GF16_inv_282_x_reg;
  wire   [8:1] Inst_GF16_inv_282_t;
  wire   [8:1] Inst_GF16_inv_282_z;
  wire   [8:1] Inst_GF16_inv_282_y;
  wire   [8:1] Inst_GF16_inv_282_x;
  wire   [4:1] Inst_Gf16_mul2_Canright1_t_reg;
  wire   [4:1] Inst_Gf16_mul2_Canright1_z_reg;
  wire   [4:1] Inst_Gf16_mul2_Canright1_y_reg;
  wire   [4:1] Inst_Gf16_mul2_Canright1_x_reg;
  wire   [4:1] Inst_Gf16_mul2_Canright1_t;
  wire   [4:1] Inst_Gf16_mul2_Canright1_z;
  wire   [4:1] Inst_Gf16_mul2_Canright1_y;
  wire   [4:1] Inst_Gf16_mul2_Canright1_x;
  wire   [4:1] Inst_Gf16_mul2_Canright2_t_reg;
  wire   [4:1] Inst_Gf16_mul2_Canright2_z_reg;
  wire   [4:1] Inst_Gf16_mul2_Canright2_y_reg;
  wire   [4:1] Inst_Gf16_mul2_Canright2_x_reg;
  wire   [4:1] Inst_Gf16_mul2_Canright2_t;
  wire   [4:1] Inst_Gf16_mul2_Canright2_z;
  wire   [4:1] Inst_Gf16_mul2_Canright2_y;
  wire   [4:1] Inst_Gf16_mul2_Canright2_x;

  DFF_X1 GEN_reg1_s_current_state_reg_0_ ( .D(dcba1[0]), .CK(clk), .Q(
        dcba1_reg1[0]), .QN() );
  DFF_X1 GEN_reg1_s_current_state_reg_1_ ( .D(dcba1[1]), .CK(clk), .Q(
        dcba1_reg1[1]), .QN() );
  DFF_X1 GEN_reg1_s_current_state_reg_2_ ( .D(dcba1[2]), .CK(clk), .Q(
        dcba1_reg1[2]), .QN() );
  DFF_X1 GEN_reg1_s_current_state_reg_3_ ( .D(dcba1[3]), .CK(clk), .Q(
        dcba1_reg1[3]), .QN() );
  DFF_X1 GEN_reg1_s_current_state_reg_4_ ( .D(dcba2[0]), .CK(clk), .Q(
        dcba2_reg1[0]), .QN() );
  DFF_X1 GEN_reg1_s_current_state_reg_5_ ( .D(dcba2[1]), .CK(clk), .Q(
        dcba2_reg1[1]), .QN() );
  DFF_X1 GEN_reg1_s_current_state_reg_6_ ( .D(dcba2[2]), .CK(clk), .Q(
        dcba2_reg1[2]), .QN() );
  DFF_X1 GEN_reg1_s_current_state_reg_7_ ( .D(dcba2[3]), .CK(clk), .Q(
        dcba2_reg1[3]), .QN() );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U51 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n47), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n46), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_z[1]) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U50 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n45), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n44), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n46)
         );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U49 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n43), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n42), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n45) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U48 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n41), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n40), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n43) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U47 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n39), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n38), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_y[1]) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U46 ( 
        .A1(hgfe1[1]), .A2(dcba1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n38) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U45 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n37), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n36), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n39) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U44 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n35), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n40), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n36) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U43 ( 
        .A1(dcba1[1]), .A2(hgfe1[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n40) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U42 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n34), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n33), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n35) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U41 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n32), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n44), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n34) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U40 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n31), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n30), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n44) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U39 ( 
        .A1(hgfe1[1]), .A2(dcba1[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n30) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U38 ( 
        .A1(dcba1[0]), .A2(hgfe1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n31) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U37 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n29), .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n28), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n32) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U36 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n41), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n27), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n28)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U35 ( 
        .A1(hgfe1[0]), .A2(dcba1[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n27) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U34 ( 
        .A1(hgfe1[0]), .A2(dcba1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n41) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U33 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n26), .A2(hgfe1[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n29) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U32 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n25), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n47), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_x[1]) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U31 ( 
        .A1(hgfe1[1]), .A2(dcba1[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n33) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U30 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n23), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n22), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n25) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U29 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n37), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n21), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n22)
         );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U28 ( 
        .A(dcba1[1]), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n20), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n21)
         );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U27 ( 
        .A1(dcba1[3]), .A2(hgfe1[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n20) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U26 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n19), .A2(hgfe1[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n23) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U25 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n18), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n17), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_t[1]) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U24 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n16), .A2(hgfe1[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n17) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U23 ( 
        .A(dcba1[3]), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n26), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n16) );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U22 ( 
        .A(dcba1[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n26) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U21 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n15), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n14), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n18)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U20 ( 
        .A1(hgfe1[0]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n13), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n14) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U19 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n19), 
        .B(dcba1[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n13) );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U18 ( 
        .A(dcba1[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n19) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U17 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n12), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n11), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n15) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U16 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n24), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n10), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n11) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U15 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n37), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n9), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n10)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U14 ( 
        .A1(dcba1[2]), .A2(hgfe1[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n9) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U13 ( 
        .A1(hgfe1[3]), .A2(dcba1[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n37) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U12 ( 
        .A1(dcba1[0]), .A2(hgfe1[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n24) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U11 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n42), 
        .B(FreshRadnom), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n12) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U10 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n8), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n7), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n42)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U9 ( 
        .A1(dcba1[3]), .A2(hgfe1[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n7) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U8 ( 
        .A1(dcba1[2]), .A2(hgfe1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n8) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U7 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n5), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n6), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n47) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U6 ( 
        .A1(hgfe1[3]), .A2(dcba1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n6) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U5 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n33), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n4), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n5)
         );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U4 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n3), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n24), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n4)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U3 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n2), 
        .A2(hgfe1[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n3) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U2 ( 
        .A(dcba1[2]), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n1), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n2)
         );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_U1 ( 
        .A(dcba1[0]), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n26), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F1_n1)
         );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U49 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n46), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n45), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_z[2]) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U48 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n44), .A2(hgfe2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n45) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U47 ( 
        .A(dcba2[0]), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n43), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n44)
         );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U46 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n42), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n41), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n46) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U45 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n40), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n39), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n41) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U44 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n38), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n37), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n39) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U43 ( 
        .A1(hgfe2[0]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n43), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n37) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U42 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n36), .A2(hgfe1[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n38) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U41 ( 
        .A(dcba2[0]), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n35), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n36) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U40 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n34), .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n33), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n40) );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U39 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n32), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n33) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U38 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n31), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n30), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n42) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U37 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n29), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n28), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n30) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U36 ( 
        .A(dcba1[1]), .B(hgfe1[1]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n28) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U35 ( 
        .A1(dcba2[3]), .A2(hgfe2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n29) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U34 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n27), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n26), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_y[2]) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U33 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n31), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n25), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n26) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U32 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n35), 
        .B(hgfe2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n31) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U31 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n24), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n23), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n27)
         );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U30 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n22), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n21), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n23)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U29 ( 
        .A1(dcba2[0]), .A2(hgfe2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n21) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U28 ( 
        .A1(hgfe2[0]), .A2(dcba2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n22) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U27 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n20), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n19), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n24) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U26 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n18), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n17), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n19) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U25 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n16), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n15), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n17)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U24 ( 
        .A1(hgfe1[1]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n43), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n15) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U23 ( 
        .A(dcba2[2]), .B(dcba2[3]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n43) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U22 ( 
        .A1(dcba1[1]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n20) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U21 ( 
        .A1(hgfe2[3]), .A2(dcba1[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n16) );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U20 ( 
        .A(dcba2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n35) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U19 ( 
        .A(hgfe2[0]), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n34)
         );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U18 ( 
        .A(dcba2[3]), .B(dcba1[1]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n25) );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U17 ( 
        .A(hgfe2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U16 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n18)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U15 ( 
        .A1(hgfe1[1]), .A2(dcba2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n12) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U14 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n32), .A2(hgfe2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n13) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U13 ( 
        .A(dcba2[0]), .B(dcba1[1]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n32) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U12 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n11), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n10), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_x[2]) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U11 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n18), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n3), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n11) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U10 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n8), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n9), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n10) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U9 ( 
        .A1(hgfe1[1]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n4), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n9)
         );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U8 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n14), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n7), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n8)
         );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U7 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n5), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n6), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n7)
         );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U6 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n35), .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n34), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n6)
         );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U5 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n25), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n16), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n5)
         );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U4 ( 
        .A(dcba2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n4) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U3 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n1), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n2), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n3)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U2 ( 
        .A1(dcba2[0]), .A2(hgfe2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n2) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_U1 ( 
        .A1(dcba2[3]), .A2(hgfe2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F2_n1) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U53 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n49), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n48), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_z[3]) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U52 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n47), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n46), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n48) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U51 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n45), .A2(hgfe2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n46) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U50 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n44), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n43), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n47) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U49 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n42), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n41), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n43) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U48 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n40), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n39), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n41) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U47 ( 
        .A(dcba2[1]), .B(hgfe2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n40) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U46 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n38), .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n37), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n42) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U45 ( 
        .A(hgfe2[0]), .B(hgfe2[3]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n38) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U44 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n36), .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n35), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n44) );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U43 ( 
        .A(hgfe2[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n36) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U42 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n49), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n34), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_y[3]) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U41 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n33), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n32), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n34) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U40 ( 
        .A1(hgfe2[3]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n31), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n32) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U39 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n30), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n29), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n33)
         );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U38 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n28), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n27), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n29) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U37 ( 
        .A1(dcba2[1]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n26), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n27) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U36 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25), .A2(hgfe2[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n28) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U35 ( 
        .A(dcba1[0]), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n37), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n25)
         );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U34 ( 
        .A1(dcba1[3]), .A2(hgfe2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n30) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U33 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n49)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U32 ( 
        .A1(hgfe2[3]), .A2(dcba1[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n23) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U31 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_x[3]) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U30 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n21) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U29 ( 
        .A(hgfe2[0]), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n37), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n19) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U28 ( 
        .A(dcba1[3]), .B(dcba1[2]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n37) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U27 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18), .A2(hgfe2[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n20) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U26 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n17), 
        .B(dcba1[3]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n18) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U25 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n16), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n15), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n22) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U24 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n14), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n13), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n15)
         );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U23 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n12), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n11), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n13)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U22 ( 
        .A1(hgfe2[3]), .A2(dcba1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n11) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U21 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n10), .A2(dcba1[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n12) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U20 ( 
        .A(hgfe2[0]), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n26), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n10) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U19 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n31), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n14)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U18 ( 
        .A1(hgfe2[0]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n45), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n24) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U17 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n17), 
        .B(dcba2[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n45) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U16 ( 
        .A1(dcba1[0]), .A2(hgfe2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n16) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U15 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n9), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n8), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_t[3]) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U14 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n31), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n39), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n8)
         );
  AND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U13 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n26), .A2(dcba1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n39) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U12 ( 
        .A1(dcba2[1]), .A2(hgfe2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n31) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U11 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n7), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n6), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n9)
         );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U10 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n5), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n4), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n6)
         );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U9 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n3), 
        .B(hgfe2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n4) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U8 ( 
        .A1(hgfe2[3]), .A2(dcba1[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n3) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U7 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n2), 
        .A2(hgfe2[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n5) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U6 ( 
        .A(dcba1[3]), .B(dcba2[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n2) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U5 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n1), 
        .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n35), .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n7) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U4 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n17), 
        .B(dcba1[2]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n35) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U3 ( 
        .A(hgfe2[0]), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n26), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n1)
         );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U2 ( 
        .A(hgfe2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n26) );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_U1 ( 
        .A(dcba1[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F3_n17) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U47 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n44), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n43), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_z[4]) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U46 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n42), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n41), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n43) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U45 ( 
        .A1(hgfe1[2]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n40), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n41) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U44 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n39), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n38), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n42)
         );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U43 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n37), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n36), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n38) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U42 ( 
        .A1(hgfe1[3]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n35), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n36) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U41 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n34), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n33), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n37)
         );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U40 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n32), .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n31), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n33) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U39 ( 
        .A(hgfe1[0]), .B(hgfe1[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n32) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U38 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n30), .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n29), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n34) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U37 ( 
        .A(hgfe1[0]), .B(hgfe1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n29) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U36 ( 
        .A(dcba2[3]), .B(dcba2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n30) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U35 ( 
        .A(dcba2[0]), .B(hgfe1[0]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n39) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U34 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n28), .A2(hgfe2[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n44) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U33 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n35), 
        .B(dcba2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n28) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U32 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n27), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n26), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_y[4]) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U31 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n25), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n24), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n26) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U30 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n23), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n22), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n24)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U29 ( 
        .A1(hgfe1[0]), .A2(dcba2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n22) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U28 ( 
        .A1(dcba2[1]), .A2(hgfe1[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n23) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U27 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n21), .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n20), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n25) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U26 ( 
        .A1(hgfe1[0]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n19), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n20) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U25 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n31), .A2(hgfe1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n21) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U24 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n18), .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n17), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n27) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U23 ( 
        .A1(hgfe2[1]), .A2(dcba2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n17) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U22 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n16), .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n15), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n18) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U21 ( 
        .A1(dcba2[3]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n35), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n15) );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U20 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n19), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n31) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U19 ( 
        .A(dcba2[0]), .B(dcba2[1]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n19) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U18 ( 
        .A1(hgfe2[1]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n14), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n16) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U17 ( 
        .A1(dcba2[3]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n35), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n14) );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U16 ( 
        .A(dcba2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n40) );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U15 ( 
        .A(dcba2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n35) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U14 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n13), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n12), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_x[4]) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U13 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n31), .A2(hgfe1[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n13) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U12 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n10), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n11), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n12) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U11 ( 
        .A1(dcba2[1]), .A2(hgfe1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n11) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U10 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n4), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n9), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n10) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U9 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n7), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n8), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n9)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U8 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n5), 
        .A2(dcba2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n8) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U7 ( 
        .A1(hgfe1[2]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n6), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n7)
         );
  INV_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U6 ( 
        .A(dcba2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n6) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U5 ( 
        .A(hgfe1[0]), .B(hgfe1[2]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n5) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U4 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n2), 
        .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n3), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n4)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U3 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n40), .A2(dcba2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n3) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U2 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n1), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n16), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n2)
         );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_U1 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n40), .A2(hgfe1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F4_n1) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U13 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n12), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n11), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_t[2]) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U12 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n10), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n9), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n11) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U11 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n8), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n7), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n9)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U10 ( 
        .A1(hgfe1[2]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n6), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n7)
         );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U9 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n5), 
        .B(dcba2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n6) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U8 ( 
        .A(dcba2[2]), .B(dcba2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n5) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U7 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n4), 
        .A2(hgfe2[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n8) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U6 ( 
        .A(dcba2[3]), .B(dcba1[1]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n4) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U5 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n3), 
        .A2(hgfe2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n10) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U4 ( 
        .A(dcba2[2]), .B(dcba2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n3) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U3 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n2), 
        .A2(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n1), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n12) );
  AND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U2 ( 
        .A1(dcba2[2]), .A2(hgfe2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n1) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_U1 ( 
        .A1(dcba1[1]), .A2(hgfe2[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F5_n2) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U15 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n34), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n33), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_t[4]) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U14 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n32), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n31), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n33)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U13 ( 
        .A1(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n30), .A2(hgfe2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n31) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U12 ( 
        .A(dcba2[3]), .B(dcba2[0]), .Z(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n30) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U11 ( 
        .A1(dcba2[2]), .A2(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n29), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n32) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U10 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n28), 
        .B(hgfe2[2]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n29) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U9 ( 
        .A(hgfe1[0]), .B(hgfe1[3]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n28) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U8 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n27), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n26), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n34) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U7 ( 
        .A1(dcba2[3]), .A2(hgfe1[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n26) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U6 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n25), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n24), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n27) );
  XNOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U5 ( 
        .A(FreshRadnom), .B(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n23), 
        .ZN(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n24) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U4 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n22), 
        .B(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n21), 
        .Z(Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n23)
         );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U3 ( 
        .A1(hgfe1[0]), .A2(dcba2[0]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n21) );
  NOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U2 ( 
        .A1(hgfe1[3]), .A2(dcba2[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n22) );
  NAND2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_U1 ( 
        .A1(hgfe1[1]), .A2(dcba2[1]), .ZN(
        Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_N_F6_n25) );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_0_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_x[1]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_x_reg[1]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_1_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_x[2]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_x_reg[2]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_2_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_x[3]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_x_reg[3]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_3_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_x[4]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_x_reg[4]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_4_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_y[1]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_y_reg[1]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_5_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_y[2]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_y_reg[2]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_6_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_y[3]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_y_reg[3]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_7_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_y[4]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_y_reg[4]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_8_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_z[1]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_z_reg[1]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_9_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_z[2]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_z_reg[2]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_10_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_z[3]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_z_reg[3]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_11_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_z[4]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_z_reg[4]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_12_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_t[1]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_t_reg[1]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_13_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_t[2]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_t_reg[2]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_14_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_t[3]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_t_reg[3]), .QN() );
  DFF_X1 Inst_Gf6_sq_scl_mul_Canright_GEN_reg_s_current_state_reg_15_ ( .D(
        Inst_Gf6_sq_scl_mul_Canright_t[4]), .CK(clk), .Q(
        Inst_Gf6_sq_scl_mul_Canright_t_reg[4]), .QN() );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L_XORInst0_U1 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_x_reg[1]), .B(
        Inst_Gf6_sq_scl_mul_Canright_x_reg[2]), .Z(sq_scl_mul_out1[1]) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U1 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_x_reg[3]), .B(
        Inst_Gf6_sq_scl_mul_Canright_x_reg[4]), .Z(sq_scl_mul_out2[1]) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U1 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_y_reg[1]), .B(
        Inst_Gf6_sq_scl_mul_Canright_y_reg[2]), .Z(sq_scl_mul_out1[2]) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U1 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_y_reg[3]), .B(
        Inst_Gf6_sq_scl_mul_Canright_y_reg[4]), .Z(sq_scl_mul_out2[2]) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U1 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_z_reg[1]), .B(
        Inst_Gf6_sq_scl_mul_Canright_z_reg[2]), .Z(sq_scl_mul_out1[3]) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U1 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_z_reg[3]), .B(
        Inst_Gf6_sq_scl_mul_Canright_z_reg[4]), .Z(sq_scl_mul_out2[3]) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U1 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_t_reg[1]), .B(
        Inst_Gf6_sq_scl_mul_Canright_t_reg[2]), .Z(sq_scl_mul_out1[4]) );
  XOR2_X1 Inst_Gf6_sq_scl_mul_Canright_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U1 ( 
        .A(Inst_Gf6_sq_scl_mul_Canright_t_reg[3]), .B(
        Inst_Gf6_sq_scl_mul_Canright_t_reg[4]), .Z(sq_scl_mul_out2[4]) );
  DFF_X1 GEN_reg2_s_current_state_reg_0_ ( .D(hgfe1[0]), .CK(clk), .Q(
        hgfe1_reg1[0]), .QN() );
  DFF_X1 GEN_reg2_s_current_state_reg_1_ ( .D(hgfe1[1]), .CK(clk), .Q(
        hgfe1_reg1[1]), .QN() );
  DFF_X1 GEN_reg2_s_current_state_reg_2_ ( .D(hgfe1[2]), .CK(clk), .Q(
        hgfe1_reg1[2]), .QN() );
  DFF_X1 GEN_reg2_s_current_state_reg_3_ ( .D(hgfe1[3]), .CK(clk), .Q(
        hgfe1_reg1[3]), .QN() );
  DFF_X1 GEN_reg2_s_current_state_reg_4_ ( .D(hgfe2[0]), .CK(clk), .Q(
        hgfe2_reg1[0]), .QN() );
  DFF_X1 GEN_reg2_s_current_state_reg_5_ ( .D(hgfe2[1]), .CK(clk), .Q(
        hgfe2_reg1[1]), .QN() );
  DFF_X1 GEN_reg2_s_current_state_reg_6_ ( .D(hgfe2[2]), .CK(clk), .Q(
        hgfe2_reg1[2]), .QN() );
  DFF_X1 GEN_reg2_s_current_state_reg_7_ ( .D(hgfe2[3]), .CK(clk), .Q(
        hgfe2_reg1[3]), .QN() );
  DFF_X1 GEN_reg3_s_current_state_reg_0_ ( .D(dcba1_reg1[0]), .CK(clk), .Q(
        dcba1_reg2[0]), .QN() );
  DFF_X1 GEN_reg3_s_current_state_reg_1_ ( .D(dcba1_reg1[1]), .CK(clk), .Q(
        dcba1_reg2[1]), .QN() );
  DFF_X1 GEN_reg3_s_current_state_reg_2_ ( .D(dcba1_reg1[2]), .CK(clk), .Q(
        dcba1_reg2[2]), .QN() );
  DFF_X1 GEN_reg3_s_current_state_reg_3_ ( .D(dcba1_reg1[3]), .CK(clk), .Q(
        dcba1_reg2[3]), .QN() );
  DFF_X1 GEN_reg3_s_current_state_reg_4_ ( .D(dcba2_reg1[0]), .CK(clk), .Q(
        dcba2_reg2[0]), .QN() );
  DFF_X1 GEN_reg3_s_current_state_reg_5_ ( .D(dcba2_reg1[1]), .CK(clk), .Q(
        dcba2_reg2[1]), .QN() );
  DFF_X1 GEN_reg3_s_current_state_reg_6_ ( .D(dcba2_reg1[2]), .CK(clk), .Q(
        dcba2_reg2[2]), .QN() );
  DFF_X1 GEN_reg3_s_current_state_reg_7_ ( .D(dcba2_reg1[3]), .CK(clk), .Q(
        dcba2_reg2[3]), .QN() );
  DFF_X1 GEN_reg4_s_current_state_reg_0_ ( .D(sq_scl_mul_out1[1]), .CK(clk), 
        .Q(sq_scl_mul_out1_reg[1]), .QN() );
  DFF_X1 GEN_reg4_s_current_state_reg_1_ ( .D(sq_scl_mul_out1[2]), .CK(clk), 
        .Q(sq_scl_mul_out1_reg[2]), .QN() );
  DFF_X1 GEN_reg4_s_current_state_reg_2_ ( .D(sq_scl_mul_out1[3]), .CK(clk), 
        .Q(sq_scl_mul_out1_reg[3]), .QN() );
  DFF_X1 GEN_reg4_s_current_state_reg_3_ ( .D(sq_scl_mul_out1[4]), .CK(clk), 
        .Q(sq_scl_mul_out1_reg[4]), .QN() );
  DFF_X1 GEN_reg4_s_current_state_reg_4_ ( .D(sq_scl_mul_out2[1]), .CK(clk), 
        .Q(sq_scl_mul_out2_reg[1]), .QN() );
  DFF_X1 GEN_reg4_s_current_state_reg_5_ ( .D(sq_scl_mul_out2[2]), .CK(clk), 
        .Q(sq_scl_mul_out2_reg[2]), .QN() );
  DFF_X1 GEN_reg4_s_current_state_reg_6_ ( .D(sq_scl_mul_out2[3]), .CK(clk), 
        .Q(sq_scl_mul_out2_reg[3]), .QN() );
  DFF_X1 GEN_reg4_s_current_state_reg_7_ ( .D(sq_scl_mul_out2[4]), .CK(clk), 
        .Q(sq_scl_mul_out2_reg[4]), .QN() );
  DFF_X1 GEN_reg5_s_current_state_reg_0_ ( .D(hgfe1_reg1[0]), .CK(clk), .Q(
        hgfe1_reg2[0]), .QN() );
  DFF_X1 GEN_reg5_s_current_state_reg_1_ ( .D(hgfe1_reg1[1]), .CK(clk), .Q(
        hgfe1_reg2[1]), .QN() );
  DFF_X1 GEN_reg5_s_current_state_reg_2_ ( .D(hgfe1_reg1[2]), .CK(clk), .Q(
        hgfe1_reg2[2]), .QN() );
  DFF_X1 GEN_reg5_s_current_state_reg_3_ ( .D(hgfe1_reg1[3]), .CK(clk), .Q(
        hgfe1_reg2[3]), .QN() );
  DFF_X1 GEN_reg5_s_current_state_reg_4_ ( .D(hgfe2_reg1[0]), .CK(clk), .Q(
        hgfe2_reg2[0]), .QN() );
  DFF_X1 GEN_reg5_s_current_state_reg_5_ ( .D(hgfe2_reg1[1]), .CK(clk), .Q(
        hgfe2_reg2[1]), .QN() );
  DFF_X1 GEN_reg5_s_current_state_reg_6_ ( .D(hgfe2_reg1[2]), .CK(clk), .Q(
        hgfe2_reg2[2]), .QN() );
  DFF_X1 GEN_reg5_s_current_state_reg_7_ ( .D(hgfe2_reg1[3]), .CK(clk), .Q(
        hgfe2_reg2[3]), .QN() );
  DFF_X1 GEN_reg6_s_current_state_reg_0_ ( .D(dcba1_reg2[0]), .CK(clk), .Q(
        dcba1_reg3[0]), .QN() );
  DFF_X1 GEN_reg6_s_current_state_reg_1_ ( .D(dcba1_reg2[1]), .CK(clk), .Q(
        dcba1_reg3[1]), .QN() );
  DFF_X1 GEN_reg6_s_current_state_reg_2_ ( .D(dcba1_reg2[2]), .CK(clk), .Q(
        dcba1_reg3[2]), .QN() );
  DFF_X1 GEN_reg6_s_current_state_reg_3_ ( .D(dcba1_reg2[3]), .CK(clk), .Q(
        dcba1_reg3[3]), .QN() );
  DFF_X1 GEN_reg6_s_current_state_reg_4_ ( .D(dcba2_reg2[0]), .CK(clk), .Q(
        dcba2_reg3[0]), .QN() );
  DFF_X1 GEN_reg6_s_current_state_reg_5_ ( .D(dcba2_reg2[1]), .CK(clk), .Q(
        dcba2_reg3[1]), .QN() );
  DFF_X1 GEN_reg6_s_current_state_reg_6_ ( .D(dcba2_reg2[2]), .CK(clk), .Q(
        dcba2_reg3[2]), .QN() );
  DFF_X1 GEN_reg6_s_current_state_reg_7_ ( .D(dcba2_reg2[3]), .CK(clk), .Q(
        dcba2_reg3[3]), .QN() );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_U4 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_n3), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_n2), .ZN(
        Inst_GF16_inv_282_x[1]) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_U3 ( .A(
        sq_scl_mul_out1_reg[2]), .B(sq_scl_mul_out1_reg[3]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_n2) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_U2 ( .A(
        sq_scl_mul_out1_reg[4]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_n1), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_n3) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_U1 ( .A1(
        sq_scl_mul_out1_reg[2]), .A2(sq_scl_mul_out1_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F1_n1) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_U4 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_n3), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_n2), .ZN(
        Inst_GF16_inv_282_x[2]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_U3 ( .A(
        sq_scl_mul_out1_reg[2]), .B(sq_scl_mul_out1_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_n2) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_U2 ( .A(
        sq_scl_mul_out2_reg[4]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_n1), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_n3) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_U1 ( .A1(
        sq_scl_mul_out2_reg[1]), .A2(sq_scl_mul_out1_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F2_n1) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U13 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n9), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n8), .ZN(
        Inst_GF16_inv_282_z[3]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U12 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n7), .A2(
        sq_scl_mul_out1_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n8) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U11 ( .A(
        sq_scl_mul_out1_reg[2]), .B(sq_scl_mul_out1_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n7) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U10 ( .A1(
        sq_scl_mul_out1_reg[1]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n6), .ZN(
        Inst_GF16_inv_282_y[3]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U9 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n5), .A2(
        sq_scl_mul_out1_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n6) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U8 ( .A(
        sq_scl_mul_out1_reg[2]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n9), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n5) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U7 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n9), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n4), .ZN(
        Inst_GF16_inv_282_x[3]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U6 ( .A(
        sq_scl_mul_out1_reg[4]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n3), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n4) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U5 ( .A1(
        sq_scl_mul_out1_reg[2]), .A2(sq_scl_mul_out1_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n3) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U4 ( .A(
        sq_scl_mul_out2_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n9) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U3 ( .A1(
        sq_scl_mul_out1_reg[2]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n2), .ZN(
        Inst_GF16_inv_282_t[3]) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U2 ( .A(
        sq_scl_mul_out1_reg[1]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n1), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n2) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_U1 ( .A1(
        sq_scl_mul_out1_reg[4]), .A2(sq_scl_mul_out2_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F3_n1) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U25 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n21), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n20), .ZN(
        Inst_GF16_inv_282_z[4]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U24 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n19), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n18), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n20) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U23 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n17), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n16), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n18) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U22 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n15), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n17), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n19) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U21 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n14), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n13), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n17) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U20 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n12), .A2(
        sq_scl_mul_out2_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n14) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U19 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n11), .B(
        sq_scl_mul_out2_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n12) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U18 ( .A1(
        sq_scl_mul_out1_reg[2]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n16), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n11) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U17 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n10), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n9), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n15) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U16 ( .A1(
        sq_scl_mul_out2_reg[1]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n8), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n21) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U15 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n7), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n6), .ZN(
        Inst_GF16_inv_282_y[4]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U14 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n5), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n13), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n6) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U13 ( .A1(
        sq_scl_mul_out2_reg[3]), .A2(sq_scl_mul_out2_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n13) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U12 ( .A1(
        sq_scl_mul_out2_reg[4]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n4), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n5) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U11 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n8), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n7) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U10 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n9), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n16), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n8) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U9 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n3), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n16), .ZN(
        Inst_GF16_inv_282_x[4]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U8 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n4), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n9), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n3) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U7 ( .A(
        sq_scl_mul_out2_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n9) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U6 ( .A1(
        sq_scl_mul_out2_reg[1]), .A2(sq_scl_mul_out1_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n4) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U5 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n2), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n10), .ZN(
        Inst_GF16_inv_282_t[4]) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U4 ( .A(
        sq_scl_mul_out1_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n10) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U3 ( .A(
        sq_scl_mul_out2_reg[1]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n1), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n2) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U2 ( .A1(
        sq_scl_mul_out2_reg[4]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n16), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n1) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_U1 ( .A(
        sq_scl_mul_out2_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F4_n16) );
  AND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_U5 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n4), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n3), .ZN(
        Inst_GF16_inv_282_x[5]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_U4 ( .A1(
        sq_scl_mul_out1_reg[3]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n2), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n3) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_U3 ( .A(
        sq_scl_mul_out2_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n2) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_U2 ( .A(
        sq_scl_mul_out2_reg[1]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n1), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n4) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_U1 ( .A1(
        sq_scl_mul_out2_reg[2]), .A2(sq_scl_mul_out1_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F5_n1) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U18 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n14), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n13), .ZN(
        Inst_GF16_inv_282_z[5]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U17 ( .A1(
        sq_scl_mul_out2_reg[2]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n12), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n13) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U16 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n11), .A2(
        sq_scl_mul_out1_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n14) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U15 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n10), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n9), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n11) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U14 ( .A1(
        sq_scl_mul_out1_reg[1]), .A2(sq_scl_mul_out1_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n9) );
  OR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U13 ( .A1(
        sq_scl_mul_out1_reg[3]), .A2(sq_scl_mul_out2_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n10) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U12 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n8), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n7), .ZN(
        Inst_GF16_inv_282_y[5]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U11 ( .A1(
        sq_scl_mul_out1_reg[1]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n12), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n7) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U10 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n6), .B(
        sq_scl_mul_out2_reg[2]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n8) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U9 ( .A1(
        sq_scl_mul_out1_reg[1]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n5), .ZN(
        Inst_GF16_inv_282_x[6]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U8 ( .A1(
        sq_scl_mul_out2_reg[2]), .A2(sq_scl_mul_out1_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n5) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U7 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n4), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n3), .ZN(
        Inst_GF16_inv_282_t[5]) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U6 ( .A1(
        sq_scl_mul_out1_reg[4]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n2), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n3) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U5 ( .A(
        sq_scl_mul_out1_reg[1]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n1), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n2) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U4 ( .A1(
        sq_scl_mul_out2_reg[2]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n6), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n1) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U3 ( .A(
        sq_scl_mul_out1_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n6) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U2 ( .A1(
        sq_scl_mul_out2_reg[2]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n12), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n4) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_U1 ( .A(
        sq_scl_mul_out1_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F6_n12) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U13 ( .A1(
        sq_scl_mul_out1_reg[4]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n9), .ZN(
        Inst_GF16_inv_282_z[7]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U12 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n8), .A2(
        sq_scl_mul_out2_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n9) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U11 ( .A(
        sq_scl_mul_out2_reg[1]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n7), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n8) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U10 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n6), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n5), .ZN(
        Inst_GF16_inv_282_y[7]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U9 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n4), .A2(
        sq_scl_mul_out1_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n5) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U8 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n7), .B(
        sq_scl_mul_out2_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n6) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U7 ( .A1(
        sq_scl_mul_out2_reg[1]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n3), .ZN(
        Inst_GF16_inv_282_x[7]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U6 ( .A1(
        sq_scl_mul_out2_reg[3]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n7), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n3) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U5 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n2), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n4), .ZN(
        Inst_GF16_inv_282_t[7]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U4 ( .A1(
        sq_scl_mul_out2_reg[1]), .A2(sq_scl_mul_out1_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n4) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U3 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n1), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n7), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n2) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U2 ( .A(
        sq_scl_mul_out2_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n7) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_U1 ( .A1(
        sq_scl_mul_out1_reg[4]), .A2(sq_scl_mul_out2_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F7_n1) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U15 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n11), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n10), .ZN(
        Inst_GF16_inv_282_z[8]) );
  OR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U14 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n9), .A2(
        sq_scl_mul_out2_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n10) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U13 ( .A(
        sq_scl_mul_out2_reg[2]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n8), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n11) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U12 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n7), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n6), .ZN(
        Inst_GF16_inv_282_y[8]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U11 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n5), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n4), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n6) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U10 ( .A1(
        sq_scl_mul_out2_reg[4]), .A2(sq_scl_mul_out1_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n5) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U9 ( .A1(
        sq_scl_mul_out2_reg[3]), .A2(sq_scl_mul_out2_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n7) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U8 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n3), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n4), .ZN(
        Inst_GF16_inv_282_x[8]) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U7 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n2), .B(
        sq_scl_mul_out1_reg[1]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n3) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U6 ( .A1(
        sq_scl_mul_out2_reg[2]), .A2(sq_scl_mul_out2_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n2) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U5 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n1), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n9), .ZN(
        Inst_GF16_inv_282_t[8]) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U4 ( .A(
        sq_scl_mul_out2_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n9) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U3 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n8), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n4), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n1) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U2 ( .A1(
        sq_scl_mul_out2_reg[2]), .A2(sq_scl_mul_out2_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n4) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_U1 ( .A(
        sq_scl_mul_out1_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F8_n8) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_U9 ( .A1(
        sq_scl_mul_out1_reg[4]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n6), .ZN(
        Inst_GF16_inv_282_z[1]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_U8 ( .A1(
        sq_scl_mul_out1_reg[3]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n5), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n6) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_U7 ( .A(
        sq_scl_mul_out1_reg[2]), .B(sq_scl_mul_out2_reg[1]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n5) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_U6 ( .A1(
        sq_scl_mul_out1_reg[4]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n4), .ZN(
        Inst_GF16_inv_282_y[1]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_U5 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n3), .A2(
        sq_scl_mul_out2_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n4) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_U4 ( .A(
        sq_scl_mul_out1_reg[2]), .B(sq_scl_mul_out1_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n3) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_U3 ( .A1(
        sq_scl_mul_out1_reg[2]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n2), .ZN(
        Inst_GF16_inv_282_t[1]) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_U2 ( .A(
        sq_scl_mul_out2_reg[1]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n1), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n2) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_U1 ( .A1(
        sq_scl_mul_out1_reg[4]), .A2(sq_scl_mul_out1_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F9_n1) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U15 ( .A1(
        sq_scl_mul_out1_reg[3]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n12), .ZN(
        Inst_GF16_inv_282_z[2]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U14 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n11), .A2(
        sq_scl_mul_out2_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n12) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U13 ( .A(
        sq_scl_mul_out1_reg[1]), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n10), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n11) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U12 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n9), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n8), .ZN(
        Inst_GF16_inv_282_y[2]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U11 ( .A1(
        sq_scl_mul_out2_reg[4]), .A2(sq_scl_mul_out1_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n8) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U10 ( .A(
        sq_scl_mul_out1_reg[3]), .B(sq_scl_mul_out1_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n9) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U9 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n7), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n6), .ZN(
        Inst_GF16_inv_282_t[2]) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U8 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n5), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n4), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n6) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U7 ( .A1(
        sq_scl_mul_out1_reg[3]), .A2(sq_scl_mul_out2_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n4) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U6 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n3), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n10), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n5) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U5 ( .A(
        sq_scl_mul_out1_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n10) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U4 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n2), .A2(
        sq_scl_mul_out2_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n7) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U3 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n1), .A2(
        sq_scl_mul_out1_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n2) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U2 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n3), .A2(
        sq_scl_mul_out1_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n1) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_U1 ( .A(
        sq_scl_mul_out1_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F10_n3) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U13 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n10), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n9), .ZN(
        Inst_GF16_inv_282_z[6]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U12 ( .A(
        sq_scl_mul_out2_reg[1]), .B(sq_scl_mul_out2_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n10) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U11 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n9), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n8), .ZN(
        Inst_GF16_inv_282_y[6]) );
  AND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U10 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n7), .A2(
        sq_scl_mul_out2_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n8) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U9 ( .A1(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n6), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n5), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n7) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U8 ( .A1(
        sq_scl_mul_out2_reg[1]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n4), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n5) );
  NAND2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U7 ( .A1(
        sq_scl_mul_out1_reg[3]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n3), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n6) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U6 ( .A(
        sq_scl_mul_out2_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n3) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U5 ( .A1(
        sq_scl_mul_out2_reg[4]), .A2(sq_scl_mul_out1_reg[3]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n9) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U4 ( .A1(
        sq_scl_mul_out2_reg[4]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n2), .ZN(
        Inst_GF16_inv_282_t[6]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U3 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n1), .B(
        sq_scl_mul_out2_reg[1]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n2) );
  NOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U2 ( .A1(
        sq_scl_mul_out1_reg[3]), .A2(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n4), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n1) );
  INV_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_U1 ( .A(
        sq_scl_mul_out2_reg[2]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_N_F11_n4) );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_0_ ( .D(
        Inst_GF16_inv_282_x[1]), .CK(clk), .Q(Inst_GF16_inv_282_x_reg[1]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_1_ ( .D(
        Inst_GF16_inv_282_x[2]), .CK(clk), .Q(Inst_GF16_inv_282_x_reg[2]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_2_ ( .D(
        Inst_GF16_inv_282_x[3]), .CK(clk), .Q(Inst_GF16_inv_282_x_reg[3]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_3_ ( .D(
        Inst_GF16_inv_282_x[4]), .CK(clk), .Q(Inst_GF16_inv_282_x_reg[4]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_4_ ( .D(
        Inst_GF16_inv_282_x[5]), .CK(clk), .Q(Inst_GF16_inv_282_x_reg[5]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_5_ ( .D(
        Inst_GF16_inv_282_x[6]), .CK(clk), .Q(Inst_GF16_inv_282_x_reg[6]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_6_ ( .D(
        Inst_GF16_inv_282_x[7]), .CK(clk), .Q(Inst_GF16_inv_282_x_reg[7]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_7_ ( .D(
        Inst_GF16_inv_282_x[8]), .CK(clk), .Q(Inst_GF16_inv_282_x_reg[8]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_8_ ( .D(
        Inst_GF16_inv_282_y[1]), .CK(clk), .Q(Inst_GF16_inv_282_y_reg[1]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_9_ ( .D(
        Inst_GF16_inv_282_y[2]), .CK(clk), .Q(Inst_GF16_inv_282_y_reg[2]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_10_ ( .D(
        Inst_GF16_inv_282_y[3]), .CK(clk), .Q(Inst_GF16_inv_282_y_reg[3]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_11_ ( .D(
        Inst_GF16_inv_282_y[4]), .CK(clk), .Q(Inst_GF16_inv_282_y_reg[4]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_12_ ( .D(
        Inst_GF16_inv_282_y[5]), .CK(clk), .Q(Inst_GF16_inv_282_y_reg[5]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_13_ ( .D(
        Inst_GF16_inv_282_y[6]), .CK(clk), .Q(Inst_GF16_inv_282_y_reg[6]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_14_ ( .D(
        Inst_GF16_inv_282_y[7]), .CK(clk), .Q(Inst_GF16_inv_282_y_reg[7]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_15_ ( .D(
        Inst_GF16_inv_282_y[8]), .CK(clk), .Q(Inst_GF16_inv_282_y_reg[8]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_16_ ( .D(
        Inst_GF16_inv_282_z[1]), .CK(clk), .Q(Inst_GF16_inv_282_z_reg[1]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_17_ ( .D(
        Inst_GF16_inv_282_z[2]), .CK(clk), .Q(Inst_GF16_inv_282_z_reg[2]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_18_ ( .D(
        Inst_GF16_inv_282_z[3]), .CK(clk), .Q(Inst_GF16_inv_282_z_reg[3]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_19_ ( .D(
        Inst_GF16_inv_282_z[4]), .CK(clk), .Q(Inst_GF16_inv_282_z_reg[4]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_20_ ( .D(
        Inst_GF16_inv_282_z[5]), .CK(clk), .Q(Inst_GF16_inv_282_z_reg[5]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_21_ ( .D(
        Inst_GF16_inv_282_z[6]), .CK(clk), .Q(Inst_GF16_inv_282_z_reg[6]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_22_ ( .D(
        Inst_GF16_inv_282_z[7]), .CK(clk), .Q(Inst_GF16_inv_282_z_reg[7]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_23_ ( .D(
        Inst_GF16_inv_282_z[8]), .CK(clk), .Q(Inst_GF16_inv_282_z_reg[8]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_24_ ( .D(
        Inst_GF16_inv_282_t[1]), .CK(clk), .Q(Inst_GF16_inv_282_t_reg[1]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_25_ ( .D(
        Inst_GF16_inv_282_t[2]), .CK(clk), .Q(Inst_GF16_inv_282_t_reg[2]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_26_ ( .D(
        Inst_GF16_inv_282_t[3]), .CK(clk), .Q(Inst_GF16_inv_282_t_reg[3]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_27_ ( .D(
        Inst_GF16_inv_282_t[4]), .CK(clk), .Q(Inst_GF16_inv_282_t_reg[4]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_28_ ( .D(
        Inst_GF16_inv_282_t[5]), .CK(clk), .Q(Inst_GF16_inv_282_t_reg[5]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_29_ ( .D(
        Inst_GF16_inv_282_t[6]), .CK(clk), .Q(Inst_GF16_inv_282_t_reg[6]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_30_ ( .D(
        Inst_GF16_inv_282_t[7]), .CK(clk), .Q(Inst_GF16_inv_282_t_reg[7]), 
        .QN() );
  DFF_X1 Inst_GF16_inv_282_GEN_reg_s_current_state_reg_31_ ( .D(
        Inst_GF16_inv_282_t[8]), .CK(clk), .Q(Inst_GF16_inv_282_t_reg[8]), 
        .QN() );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U3 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n6), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n5), .ZN(
        GF16_inv_out1[0]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U2 ( .A(
        Inst_GF16_inv_282_x_reg[3]), .B(Inst_GF16_inv_282_x_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n5) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U1 ( .A(
        Inst_GF16_inv_282_x_reg[1]), .B(Inst_GF16_inv_282_x_reg[2]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_n6) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U3 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n6), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n5), .ZN(
        GF16_inv_out2[0]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U2 ( .A(
        Inst_GF16_inv_282_x_reg[7]), .B(Inst_GF16_inv_282_x_reg[8]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n5) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U1 ( .A(
        Inst_GF16_inv_282_x_reg[5]), .B(Inst_GF16_inv_282_x_reg[6]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_n6) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U3 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n6), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n5), .ZN(
        GF16_inv_out1[1]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U2 ( .A(
        Inst_GF16_inv_282_y_reg[3]), .B(Inst_GF16_inv_282_y_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n5) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U1 ( .A(
        Inst_GF16_inv_282_y_reg[1]), .B(Inst_GF16_inv_282_y_reg[2]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_n6) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U3 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n6), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n5), .ZN(
        GF16_inv_out2[1]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U2 ( .A(
        Inst_GF16_inv_282_y_reg[7]), .B(Inst_GF16_inv_282_y_reg[8]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n5) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U1 ( .A(
        Inst_GF16_inv_282_y_reg[5]), .B(Inst_GF16_inv_282_y_reg[6]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_n6) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U3 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n6), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n5), .ZN(
        GF16_inv_out1[2]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U2 ( .A(
        Inst_GF16_inv_282_z_reg[3]), .B(Inst_GF16_inv_282_z_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n5) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U1 ( .A(
        Inst_GF16_inv_282_z_reg[1]), .B(Inst_GF16_inv_282_z_reg[2]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_n6) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U3 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n6), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n5), .ZN(
        GF16_inv_out2[2]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U2 ( .A(
        Inst_GF16_inv_282_z_reg[7]), .B(Inst_GF16_inv_282_z_reg[8]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n5) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U1 ( .A(
        Inst_GF16_inv_282_z_reg[5]), .B(Inst_GF16_inv_282_z_reg[6]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_n6) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U3 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n6), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n5), .ZN(
        GF16_inv_out1[3]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U2 ( .A(
        Inst_GF16_inv_282_t_reg[3]), .B(Inst_GF16_inv_282_t_reg[4]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n5) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U1 ( .A(
        Inst_GF16_inv_282_t_reg[1]), .B(Inst_GF16_inv_282_t_reg[2]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_n6) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_U3 ( .A(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n6), .B(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n5), .ZN(
        GF16_inv_out2[3]) );
  XNOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_U2 ( .A(
        Inst_GF16_inv_282_t_reg[7]), .B(Inst_GF16_inv_282_t_reg[8]), .ZN(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n5) );
  XOR2_X1 Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_U1 ( .A(
        Inst_GF16_inv_282_t_reg[5]), .B(Inst_GF16_inv_282_t_reg[6]), .Z(
        Inst_GF16_inv_282_Inst_Gf6_sq_scl_mul_Canright_L_XORInst8_n6) );
  DFF_X1 GEN_reg7_s_current_state_reg_0_ ( .D(hgfe1_reg2[0]), .CK(clk), .Q(
        hgfe1_reg3[0]), .QN() );
  DFF_X1 GEN_reg7_s_current_state_reg_1_ ( .D(hgfe1_reg2[1]), .CK(clk), .Q(
        hgfe1_reg3[1]), .QN() );
  DFF_X1 GEN_reg7_s_current_state_reg_2_ ( .D(hgfe1_reg2[2]), .CK(clk), .Q(
        hgfe1_reg3[2]), .QN() );
  DFF_X1 GEN_reg7_s_current_state_reg_3_ ( .D(hgfe1_reg2[3]), .CK(clk), .Q(
        hgfe1_reg3[3]), .QN() );
  DFF_X1 GEN_reg7_s_current_state_reg_4_ ( .D(hgfe2_reg2[0]), .CK(clk), .Q(
        hgfe2_reg3[0]), .QN() );
  DFF_X1 GEN_reg7_s_current_state_reg_5_ ( .D(hgfe2_reg2[1]), .CK(clk), .Q(
        hgfe2_reg3[1]), .QN() );
  DFF_X1 GEN_reg7_s_current_state_reg_6_ ( .D(hgfe2_reg2[2]), .CK(clk), .Q(
        hgfe2_reg3[2]), .QN() );
  DFF_X1 GEN_reg7_s_current_state_reg_7_ ( .D(hgfe2_reg2[3]), .CK(clk), .Q(
        hgfe2_reg3[3]), .QN() );
  DFF_X1 GEN_reg8_s_current_state_reg_0_ ( .D(dcba1_reg3[0]), .CK(clk), .Q(
        dcba1_reg4[0]), .QN() );
  DFF_X1 GEN_reg8_s_current_state_reg_1_ ( .D(dcba1_reg3[1]), .CK(clk), .Q(
        dcba1_reg4[1]), .QN() );
  DFF_X1 GEN_reg8_s_current_state_reg_2_ ( .D(dcba1_reg3[2]), .CK(clk), .Q(
        dcba1_reg4[2]), .QN() );
  DFF_X1 GEN_reg8_s_current_state_reg_3_ ( .D(dcba1_reg3[3]), .CK(clk), .Q(
        dcba1_reg4[3]), .QN() );
  DFF_X1 GEN_reg8_s_current_state_reg_4_ ( .D(dcba2_reg3[0]), .CK(clk), .Q(
        dcba2_reg4[0]), .QN() );
  DFF_X1 GEN_reg8_s_current_state_reg_5_ ( .D(dcba2_reg3[1]), .CK(clk), .Q(
        dcba2_reg4[1]), .QN() );
  DFF_X1 GEN_reg8_s_current_state_reg_6_ ( .D(dcba2_reg3[2]), .CK(clk), .Q(
        dcba2_reg4[2]), .QN() );
  DFF_X1 GEN_reg8_s_current_state_reg_7_ ( .D(dcba2_reg3[3]), .CK(clk), .Q(
        dcba2_reg4[3]), .QN() );
  DFF_X1 GEN_reg9_s_current_state_reg_0_ ( .D(GF16_inv_out1[0]), .CK(clk), .Q(
        GF16_inv_out1_reg[0]), .QN() );
  DFF_X1 GEN_reg9_s_current_state_reg_1_ ( .D(GF16_inv_out1[1]), .CK(clk), .Q(
        GF16_inv_out1_reg[1]), .QN() );
  DFF_X1 GEN_reg9_s_current_state_reg_2_ ( .D(GF16_inv_out1[2]), .CK(clk), .Q(
        GF16_inv_out1_reg[2]), .QN() );
  DFF_X1 GEN_reg9_s_current_state_reg_3_ ( .D(GF16_inv_out1[3]), .CK(clk), .Q(
        GF16_inv_out1_reg[3]), .QN() );
  DFF_X1 GEN_reg9_s_current_state_reg_4_ ( .D(GF16_inv_out2[0]), .CK(clk), .Q(
        GF16_inv_out2_reg[0]), .QN() );
  DFF_X1 GEN_reg9_s_current_state_reg_5_ ( .D(GF16_inv_out2[1]), .CK(clk), .Q(
        GF16_inv_out2_reg[1]), .QN() );
  DFF_X1 GEN_reg9_s_current_state_reg_6_ ( .D(GF16_inv_out2[2]), .CK(clk), .Q(
        GF16_inv_out2_reg[2]), .QN() );
  DFF_X1 GEN_reg9_s_current_state_reg_7_ ( .D(GF16_inv_out2[3]), .CK(clk), .Q(
        GF16_inv_out2_reg[3]), .QN() );
  DFF_X1 GEN_reg10_s_current_state_reg_0_ ( .D(hgfe1_reg3[0]), .CK(clk), .Q(
        hgfe1_reg4[0]), .QN() );
  DFF_X1 GEN_reg10_s_current_state_reg_1_ ( .D(hgfe1_reg3[1]), .CK(clk), .Q(
        hgfe1_reg4[1]), .QN() );
  DFF_X1 GEN_reg10_s_current_state_reg_2_ ( .D(hgfe1_reg3[2]), .CK(clk), .Q(
        hgfe1_reg4[2]), .QN() );
  DFF_X1 GEN_reg10_s_current_state_reg_3_ ( .D(hgfe1_reg3[3]), .CK(clk), .Q(
        hgfe1_reg4[3]), .QN() );
  DFF_X1 GEN_reg10_s_current_state_reg_4_ ( .D(hgfe2_reg3[0]), .CK(clk), .Q(
        hgfe2_reg4[0]), .QN() );
  DFF_X1 GEN_reg10_s_current_state_reg_5_ ( .D(hgfe2_reg3[1]), .CK(clk), .Q(
        hgfe2_reg4[1]), .QN() );
  DFF_X1 GEN_reg10_s_current_state_reg_6_ ( .D(hgfe2_reg3[2]), .CK(clk), .Q(
        hgfe2_reg4[2]), .QN() );
  DFF_X1 GEN_reg10_s_current_state_reg_7_ ( .D(hgfe2_reg3[3]), .CK(clk), .Q(
        hgfe2_reg4[3]), .QN() );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U43 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126), .Z(
        Inst_Gf16_mul2_Canright1_z[1]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U42 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U41 ( 
        .A1(dcba1_reg4[3]), .A2(GF16_inv_out1_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U40 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U39 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U38 ( 
        .A1(GF16_inv_out1_reg[2]), .A2(dcba1_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U37 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U36 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116), 
        .ZN(Inst_Gf16_mul2_Canright1_y[1]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U35 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U34 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U33 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U32 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U31 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108), 
        .B(dcba1_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U30 ( 
        .A1(dcba1_reg4[3]), .A2(GF16_inv_out1_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U29 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106), 
        .ZN(Inst_Gf16_mul2_Canright1_x[1]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U28 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U27 ( 
        .A1(dcba1_reg4[0]), .A2(GF16_inv_out1_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U26 ( 
        .A(dcba1_reg4[3]), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U25 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U24 ( 
        .A1(GF16_inv_out1_reg[3]), .A2(dcba1_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U23 ( 
        .A1(GF16_inv_out1_reg[2]), .A2(dcba1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U22 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U21 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U20 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U19 ( 
        .A1(GF16_inv_out1_reg[0]), .A2(dcba1_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U18 ( 
        .A1(GF16_inv_out1_reg[1]), .A2(dcba1_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U17 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101), 
        .ZN(Inst_Gf16_mul2_Canright1_t[1]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U16 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U15 ( 
        .A1(GF16_inv_out1_reg[1]), .A2(dcba1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U14 ( 
        .A1(GF16_inv_out1_reg[1]), .A2(dcba1_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U13 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U12 ( .A(
        dcba1_reg4[0]), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U11 ( 
        .A1(dcba1_reg4[1]), .A2(GF16_inv_out1_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U10 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U9 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91), 
        .A2(GF16_inv_out1_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U8 ( .A(
        dcba1_reg4[1]), .B(dcba1_reg4[2]), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U7 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U6 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n90), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U5 ( 
        .A1(dcba1_reg4[2]), .A2(GF16_inv_out1_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n90) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U4 ( 
        .A1(dcba1_reg4[3]), .A2(GF16_inv_out1_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U3 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n89), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U2 ( 
        .A1(GF16_inv_out1_reg[0]), .A2(dcba1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n89) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_U1 ( 
        .A1(dcba1_reg4[0]), .A2(GF16_inv_out1_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U47 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136), 
        .ZN(Inst_Gf16_mul2_Canright1_y[2]) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U46 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U45 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U44 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132), 
        .B(dcba1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U43 ( 
        .A1(dcba1_reg4[3]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U42 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131), 
        .A2(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U41 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n141), 
        .A2(GF16_inv_out2_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131) );
  INV_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U40 ( .A(
        dcba1_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n141) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U39 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128), 
        .ZN(Inst_Gf16_mul2_Canright1_x[2]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U38 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U37 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U36 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U35 ( 
        .A1(GF16_inv_out2_reg[3]), .A2(dcba1_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U34 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n142), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U33 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n142) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U32 ( 
        .A1(dcba1_reg4[0]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U31 ( 
        .A1(dcba1_reg4[0]), .A2(GF16_inv_out2_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U30 ( 
        .A(GF16_inv_out2_reg[0]), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n140), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U29 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(dcba1_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n140) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U28 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118), 
        .ZN(Inst_Gf16_mul2_Canright1_t[2]) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U27 ( 
        .A1(dcba1_reg4[1]), .A2(GF16_inv_out2_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U26 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U25 ( 
        .A1(GF16_inv_out2_reg[3]), .A2(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116) );
  INV_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U24 ( .A(
        dcba1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U23 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U22 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U21 ( 
        .A(dcba1_reg4[1]), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U20 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n143), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U19 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n143) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U18 ( .A(
        dcba1_reg4[3]), .B(dcba1_reg4[0]), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U17 ( 
        .A1(GF16_inv_out2_reg[2]), .A2(dcba1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U16 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U15 ( 
        .A1(dcba1_reg4[1]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U14 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(dcba1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U13 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115)
         );
  NOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U12 ( 
        .A1(GF16_inv_out2_reg[2]), .A2(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134) );
  INV_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U11 ( .A(
        dcba1_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U10 ( 
        .A1(dcba1_reg4[2]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U9 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108), .ZN(
        Inst_Gf16_mul2_Canright1_z[2]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U8 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U7 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U6 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n140), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U5 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104), 
        .A2(GF16_inv_out2_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U4 ( .A(
        dcba1_reg4[3]), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n141), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U3 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102), 
        .A2(GF16_inv_out2_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U2 ( .A(
        dcba1_reg4[3]), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_U1 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n143), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n142), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U46 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n152), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n151), 
        .ZN(Inst_Gf16_mul2_Canright1_z[3]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U45 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n150), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n149), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n151)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U44 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n148), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n147), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n150)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U43 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n146), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n145), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n148)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U42 ( 
        .A1(dcba2_reg4[0]), .A2(GF16_inv_out1_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n145) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U41 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n144), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n143), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n146)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U40 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n142), 
        .A2(dcba2_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n152) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U39 ( .A(
        GF16_inv_out1_reg[0]), .B(GF16_inv_out1_reg[3]), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n142) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U38 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n141), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n140), 
        .ZN(Inst_Gf16_mul2_Canright1_y[3]) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U37 ( 
        .A1(GF16_inv_out1_reg[0]), .A2(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n140) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U36 ( .A(
        dcba2_reg4[3]), .B(dcba2_reg4[1]), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U35 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n141)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U34 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U33 ( 
        .A1(GF16_inv_out1_reg[3]), .A2(dcba2_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U32 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n143), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U31 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133), 
        .B(dcba2_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n143) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U30 ( 
        .A1(dcba2_reg4[3]), .A2(GF16_inv_out1_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U29 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131), 
        .ZN(Inst_Gf16_mul2_Canright1_x[3]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U28 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U27 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n144), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U26 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n144)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U25 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U24 ( 
        .A1(GF16_inv_out1_reg[1]), .A2(dcba2_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U23 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123), 
        .A2(GF16_inv_out1_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U22 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122), 
        .A2(dcba2_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U21 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121), 
        .B(GF16_inv_out1_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U20 ( 
        .A(dcba2_reg4[3]), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n149), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U19 ( 
        .A1(dcba2_reg4[0]), .A2(GF16_inv_out1_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n149) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U18 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120), 
        .A2(GF16_inv_out1_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U17 ( .A(
        dcba2_reg4[1]), .B(dcba2_reg4[0]), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U16 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118), 
        .ZN(Inst_Gf16_mul2_Canright1_t[3]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U15 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U14 ( 
        .A1(dcba2_reg4[3]), .A2(GF16_inv_out1_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U13 ( 
        .A(dcba2_reg4[0]), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U12 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U11 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n147), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U10 ( 
        .A1(GF16_inv_out1_reg[1]), .A2(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U9 ( .A(
        dcba2_reg4[2]), .B(dcba2_reg4[0]), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U8 ( 
        .A1(dcba2_reg4[2]), .A2(GF16_inv_out1_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n147) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U7 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113), 
        .A2(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U6 ( 
        .A1(GF16_inv_out1_reg[2]), .A2(dcba2_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U5 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121), 
        .A2(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U4 ( .A(
        dcba2_reg4[2]), .B(dcba2_reg4[3]), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134) );
  INV_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U3 ( .A(
        GF16_inv_out1_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U2 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111), 
        .A2(GF16_inv_out1_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_U1 ( .A(
        dcba2_reg4[2]), .B(dcba2_reg4[1]), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U46 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n140), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139), 
        .ZN(Inst_Gf16_mul2_Canright1_z[4]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U45 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U44 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U43 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U42 ( 
        .A1(dcba2_reg4[2]), .A2(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133) );
  NOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U41 ( 
        .A1(dcba2_reg4[3]), .A2(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U40 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n140)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U39 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U38 ( 
        .A1(GF16_inv_out2_reg[2]), .A2(dcba2_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U37 ( 
        .A1(GF16_inv_out2_reg[3]), .A2(dcba2_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U36 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125), 
        .ZN(Inst_Gf16_mul2_Canright1_y[4]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U35 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U34 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U33 ( 
        .A1(GF16_inv_out2_reg[0]), .A2(dcba2_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137) );
  NOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U32 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(dcba2_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U31 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120), 
        .ZN(Inst_Gf16_mul2_Canright1_x[4]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U30 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U29 ( 
        .A1(dcba2_reg4[1]), .A2(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118) );
  INV_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U28 ( .A(
        GF16_inv_out2_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U27 ( .A(
        GF16_inv_out2_reg[0]), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U26 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U25 ( 
        .A1(GF16_inv_out2_reg[0]), .A2(dcba2_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U24 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U23 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U22 ( 
        .A1(dcba2_reg4[1]), .A2(GF16_inv_out2_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U21 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U20 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U19 ( 
        .A1(GF16_inv_out2_reg[3]), .A2(dcba2_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U18 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108), 
        .ZN(Inst_Gf16_mul2_Canright1_t[4]) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U17 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U16 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U15 ( 
        .A1(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131), 
        .A2(dcba2_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105) );
  INV_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U14 ( .A(
        GF16_inv_out2_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U13 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U12 ( 
        .A(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103), 
        .B(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102), 
        .ZN(Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U11 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U10 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100), .Z(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U9 ( 
        .A1(dcba2_reg4[3]), .A2(GF16_inv_out2_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U8 ( 
        .A1(dcba2_reg4[1]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101) );
  XNOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U7 ( .A(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135), .B(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U6 ( 
        .A1(dcba2_reg4[2]), .A2(GF16_inv_out2_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U5 ( 
        .A1(dcba2_reg4[0]), .A2(GF16_inv_out2_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135) );
  NOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U4 ( .A1(
        dcba2_reg4[2]), .A2(GF16_inv_out2_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U3 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(dcba2_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U2 ( 
        .A1(dcba2_reg4[2]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115) );
  NAND2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_U1 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(dcba2_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113) );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_0_ ( .D(
        Inst_Gf16_mul2_Canright1_x[1]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_x_reg[1]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_1_ ( .D(
        Inst_Gf16_mul2_Canright1_x[2]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_x_reg[2]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_2_ ( .D(
        Inst_Gf16_mul2_Canright1_x[3]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_x_reg[3]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_3_ ( .D(
        Inst_Gf16_mul2_Canright1_x[4]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_x_reg[4]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_4_ ( .D(
        Inst_Gf16_mul2_Canright1_y[1]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_y_reg[1]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_5_ ( .D(
        Inst_Gf16_mul2_Canright1_y[2]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_y_reg[2]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_6_ ( .D(
        Inst_Gf16_mul2_Canright1_y[3]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_y_reg[3]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_7_ ( .D(
        Inst_Gf16_mul2_Canright1_y[4]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_y_reg[4]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_8_ ( .D(
        Inst_Gf16_mul2_Canright1_z[1]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_z_reg[1]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_9_ ( .D(
        Inst_Gf16_mul2_Canright1_z[2]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_z_reg[2]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_10_ ( .D(
        Inst_Gf16_mul2_Canright1_z[3]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_z_reg[3]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_11_ ( .D(
        Inst_Gf16_mul2_Canright1_z[4]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_z_reg[4]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_12_ ( .D(
        Inst_Gf16_mul2_Canright1_t[1]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_t_reg[1]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_13_ ( .D(
        Inst_Gf16_mul2_Canright1_t[2]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_t_reg[2]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_14_ ( .D(
        Inst_Gf16_mul2_Canright1_t[3]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_t_reg[3]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright1_GEN_reg_s_current_state_reg_15_ ( .D(
        Inst_Gf16_mul2_Canright1_t[4]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright1_t_reg[4]), .QN() );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst0_U1 ( 
        .A(Inst_Gf16_mul2_Canright1_x_reg[1]), .B(
        Inst_Gf16_mul2_Canright1_x_reg[2]), .Z(hgfe1_out[0]) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U1 ( 
        .A(Inst_Gf16_mul2_Canright1_x_reg[3]), .B(
        Inst_Gf16_mul2_Canright1_x_reg[4]), .Z(hgfe2_out[0]) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U1 ( 
        .A(Inst_Gf16_mul2_Canright1_y_reg[1]), .B(
        Inst_Gf16_mul2_Canright1_y_reg[2]), .Z(hgfe1_out[1]) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U1 ( 
        .A(Inst_Gf16_mul2_Canright1_y_reg[3]), .B(
        Inst_Gf16_mul2_Canright1_y_reg[4]), .Z(hgfe2_out[1]) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U1 ( 
        .A(Inst_Gf16_mul2_Canright1_z_reg[1]), .B(
        Inst_Gf16_mul2_Canright1_z_reg[2]), .Z(hgfe1_out[2]) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U1 ( 
        .A(Inst_Gf16_mul2_Canright1_z_reg[3]), .B(
        Inst_Gf16_mul2_Canright1_z_reg[4]), .Z(hgfe2_out[2]) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U1 ( 
        .A(Inst_Gf16_mul2_Canright1_t_reg[1]), .B(
        Inst_Gf16_mul2_Canright1_t_reg[2]), .Z(hgfe1_out[3]) );
  XOR2_X1 Inst_Gf16_mul2_Canright1_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U1 ( 
        .A(Inst_Gf16_mul2_Canright1_t_reg[3]), .B(
        Inst_Gf16_mul2_Canright1_t_reg[4]), .Z(hgfe2_out[3]) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U43 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126), .Z(
        Inst_Gf16_mul2_Canright2_z[1]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U42 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n126)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U41 ( 
        .A1(hgfe1_reg4[3]), .A2(GF16_inv_out1_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n124) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U40 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n125)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U39 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n122)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U38 ( 
        .A1(GF16_inv_out1_reg[2]), .A2(hgfe1_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n120) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U37 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n121) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U36 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116), 
        .ZN(Inst_Gf16_mul2_Canright2_y[1]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U35 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n117)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U34 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n115)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U33 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n113)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U32 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n111)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U31 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108), 
        .B(hgfe1_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n118) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U30 ( 
        .A1(hgfe1_reg4[3]), .A2(GF16_inv_out1_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n108) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U29 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106), 
        .ZN(Inst_Gf16_mul2_Canright2_x[1]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U28 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n106)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U27 ( 
        .A1(hgfe1_reg4[0]), .A2(GF16_inv_out1_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n110) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U26 ( 
        .A(hgfe1_reg4[3]), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n105) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U25 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n104) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U24 ( 
        .A1(GF16_inv_out1_reg[3]), .A2(hgfe1_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n102) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U23 ( 
        .A1(GF16_inv_out1_reg[2]), .A2(hgfe1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n103) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U22 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n107)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U21 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n119)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U20 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n99) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U19 ( 
        .A1(GF16_inv_out1_reg[0]), .A2(hgfe1_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n97) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U18 ( 
        .A1(GF16_inv_out1_reg[1]), .A2(hgfe1_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n98) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U17 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101), 
        .ZN(Inst_Gf16_mul2_Canright2_t[1]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U16 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n101)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U15 ( 
        .A1(GF16_inv_out1_reg[1]), .A2(hgfe1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n109) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U14 ( 
        .A1(GF16_inv_out1_reg[1]), .A2(hgfe1_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n123) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U13 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n96) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U12 ( .A(
        hgfe1_reg4[0]), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n116) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U11 ( 
        .A1(hgfe1_reg4[1]), .A2(GF16_inv_out1_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n94) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U10 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n95) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U9 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91), 
        .A2(GF16_inv_out1_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n92) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U8 ( .A(
        hgfe1_reg4[1]), .B(hgfe1_reg4[2]), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n91) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U7 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n93) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U6 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n90), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n127) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U5 ( 
        .A1(hgfe1_reg4[2]), .A2(GF16_inv_out1_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n90) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U4 ( 
        .A1(hgfe1_reg4[3]), .A2(GF16_inv_out1_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n114) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U3 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n89), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n100) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U2 ( 
        .A1(GF16_inv_out1_reg[0]), .A2(hgfe1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n89) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_U1 ( 
        .A1(hgfe1_reg4[0]), .A2(GF16_inv_out1_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F1_n112) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U47 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136), 
        .ZN(Inst_Gf16_mul2_Canright2_y[2]) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U46 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n136) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U45 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n137)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U44 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132), 
        .B(hgfe1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U43 ( 
        .A1(hgfe1_reg4[3]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n132) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U42 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131), 
        .A2(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n133)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U41 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n141), 
        .A2(GF16_inv_out2_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n131) );
  INV_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U40 ( .A(
        hgfe1_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n141) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U39 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128), 
        .ZN(Inst_Gf16_mul2_Canright2_x[2]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U38 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n128)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U37 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n127) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U36 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n126)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U35 ( 
        .A1(GF16_inv_out2_reg[3]), .A2(hgfe1_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n123) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U34 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n142), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n124) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U33 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n142) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U32 ( 
        .A1(hgfe1_reg4[0]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n120) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U31 ( 
        .A1(hgfe1_reg4[0]), .A2(GF16_inv_out2_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n130) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U30 ( 
        .A(GF16_inv_out2_reg[0]), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n140), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n129) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U29 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(hgfe1_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n140) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U28 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118), 
        .ZN(Inst_Gf16_mul2_Canright2_t[2]) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U27 ( 
        .A1(hgfe1_reg4[1]), .A2(GF16_inv_out2_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n118) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U26 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n119)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U25 ( 
        .A1(GF16_inv_out2_reg[3]), .A2(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n116) );
  INV_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U24 ( .A(
        hgfe1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U23 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n117)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U22 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n114)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U21 ( 
        .A(hgfe1_reg4[1]), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n122) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U20 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n143), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n113)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U19 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n143) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U18 ( .A(
        hgfe1_reg4[3]), .B(hgfe1_reg4[0]), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n111) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U17 ( 
        .A1(GF16_inv_out2_reg[2]), .A2(hgfe1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n112) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U16 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n135) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U15 ( 
        .A1(hgfe1_reg4[1]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n110) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U14 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(hgfe1_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n125) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U13 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n115)
         );
  NOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U12 ( 
        .A1(GF16_inv_out2_reg[2]), .A2(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n134) );
  INV_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U11 ( .A(
        hgfe1_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n109) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U10 ( 
        .A1(hgfe1_reg4[2]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n121) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U9 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107), .ZN(
        Inst_Gf16_mul2_Canright2_z[2]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U8 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n143), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n142), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n108) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U7 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n107) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U6 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105), 
        .A2(GF16_inv_out2_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n106) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U5 ( .A(
        hgfe1_reg4[3]), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n138), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n105) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U4 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n104) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U3 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102), 
        .A2(GF16_inv_out2_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n103) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U2 ( .A(
        hgfe1_reg4[3]), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n141), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n102) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_U1 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n140), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n139), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F2_n101) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U46 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n152), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n151), 
        .ZN(Inst_Gf16_mul2_Canright2_z[3]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U45 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n150), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n149), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n151)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U44 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n148), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n147), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n150)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U43 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n146), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n145), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n148)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U42 ( 
        .A1(hgfe2_reg4[0]), .A2(GF16_inv_out1_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n145) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U41 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n144), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n143), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n146)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U40 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n142), 
        .A2(hgfe2_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n152) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U39 ( .A(
        GF16_inv_out1_reg[0]), .B(GF16_inv_out1_reg[3]), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n142) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U38 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n141), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n140), 
        .ZN(Inst_Gf16_mul2_Canright2_y[3]) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U37 ( 
        .A1(GF16_inv_out1_reg[0]), .A2(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n140) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U36 ( .A(
        hgfe2_reg4[3]), .B(hgfe2_reg4[1]), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n139) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U35 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n141)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U34 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n137)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U33 ( 
        .A1(GF16_inv_out1_reg[3]), .A2(hgfe2_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n135) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U32 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n143), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n136) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U31 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133), 
        .B(hgfe2_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n143) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U30 ( 
        .A1(hgfe2_reg4[3]), .A2(GF16_inv_out1_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n133) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U29 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131), 
        .ZN(Inst_Gf16_mul2_Canright2_x[3]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U28 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n131)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U27 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n144), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n129)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U26 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n144)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U25 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n126)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U24 ( 
        .A1(GF16_inv_out1_reg[1]), .A2(hgfe2_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n124) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U23 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123), 
        .A2(GF16_inv_out1_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n125) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U22 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122), 
        .A2(hgfe2_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n128) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U21 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121), 
        .B(GF16_inv_out1_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n122) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U20 ( 
        .A(hgfe2_reg4[3]), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n149), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n130) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U19 ( 
        .A1(hgfe2_reg4[0]), .A2(GF16_inv_out1_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n149) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U18 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120), 
        .A2(GF16_inv_out1_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n132) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U17 ( .A(
        hgfe2_reg4[1]), .B(hgfe2_reg4[0]), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n120) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U16 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118), 
        .ZN(Inst_Gf16_mul2_Canright2_t[3]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U15 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n118)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U14 ( 
        .A1(hgfe2_reg4[3]), .A2(GF16_inv_out1_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n127) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U13 ( 
        .A(hgfe2_reg4[0]), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n117) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U12 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n116)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U11 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n147), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n114) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U10 ( 
        .A1(GF16_inv_out1_reg[1]), .A2(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n138) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U9 ( .A(
        hgfe2_reg4[2]), .B(hgfe2_reg4[0]), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n123) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U8 ( 
        .A1(hgfe2_reg4[2]), .A2(GF16_inv_out1_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n147) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U7 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113), 
        .A2(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n115)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U6 ( 
        .A1(GF16_inv_out1_reg[2]), .A2(hgfe2_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n112) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U5 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121), 
        .A2(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n113)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U4 ( .A(
        hgfe2_reg4[2]), .B(hgfe2_reg4[3]), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n134) );
  INV_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U3 ( .A(
        GF16_inv_out1_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n121) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U2 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111), 
        .A2(GF16_inv_out1_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n119) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_U1 ( .A(
        hgfe2_reg4[2]), .B(hgfe2_reg4[1]), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F3_n111) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U46 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n140), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139), 
        .ZN(Inst_Gf16_mul2_Canright2_z[4]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U45 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n139)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U44 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n138)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U43 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n136)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U42 ( 
        .A1(hgfe2_reg4[2]), .A2(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n133) );
  NOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U41 ( 
        .A1(hgfe2_reg4[3]), .A2(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n134) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U40 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n140)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U39 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n129) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U38 ( 
        .A1(GF16_inv_out2_reg[2]), .A2(hgfe2_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n127) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U37 ( 
        .A1(GF16_inv_out2_reg[3]), .A2(hgfe2_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n128) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U36 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125), 
        .ZN(Inst_Gf16_mul2_Canright2_y[4]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U35 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n125)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U34 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n124)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U33 ( 
        .A1(GF16_inv_out2_reg[0]), .A2(hgfe2_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n137) );
  NOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U32 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(hgfe2_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n122) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U31 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120), 
        .ZN(Inst_Gf16_mul2_Canright2_x[4]) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U30 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n120)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U29 ( 
        .A1(hgfe2_reg4[1]), .A2(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n118) );
  INV_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U28 ( .A(
        GF16_inv_out2_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n132) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U27 ( .A(
        GF16_inv_out2_reg[0]), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n119) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U26 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n130)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U25 ( 
        .A1(GF16_inv_out2_reg[0]), .A2(hgfe2_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n116) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U24 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n117)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U23 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n114) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U22 ( 
        .A1(hgfe2_reg4[1]), .A2(GF16_inv_out2_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n112) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U21 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n121)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U20 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n123)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U19 ( 
        .A1(GF16_inv_out2_reg[3]), .A2(hgfe2_reg4[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n110) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U18 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108), 
        .ZN(Inst_Gf16_mul2_Canright2_t[4]) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U17 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n108) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U16 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n107)
         );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U15 ( 
        .A1(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131), 
        .A2(hgfe2_reg4[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n105) );
  INV_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U14 ( .A(
        GF16_inv_out2_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n131) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U13 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n106)
         );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U12 ( 
        .A(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103), 
        .B(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102), 
        .ZN(Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n104)
         );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U11 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n102) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U10 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100), .Z(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n126) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U9 ( 
        .A1(hgfe2_reg4[3]), .A2(GF16_inv_out2_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n100) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U8 ( 
        .A1(hgfe2_reg4[1]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n101) );
  XNOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U7 ( .A(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135), .B(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n111) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U6 ( 
        .A1(hgfe2_reg4[2]), .A2(GF16_inv_out2_reg[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n99) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U5 ( 
        .A1(hgfe2_reg4[0]), .A2(GF16_inv_out2_reg[1]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n135) );
  NOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U4 ( .A1(
        hgfe2_reg4[2]), .A2(GF16_inv_out2_reg[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n103) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U3 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(hgfe2_reg4[2]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n109) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U2 ( 
        .A1(hgfe2_reg4[2]), .A2(GF16_inv_out2_reg[0]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n115) );
  NAND2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_U1 ( 
        .A1(GF16_inv_out2_reg[1]), .A2(hgfe2_reg4[3]), .ZN(
        Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_N_F4_n113) );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_0_ ( .D(
        Inst_Gf16_mul2_Canright2_x[1]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_x_reg[1]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_1_ ( .D(
        Inst_Gf16_mul2_Canright2_x[2]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_x_reg[2]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_2_ ( .D(
        Inst_Gf16_mul2_Canright2_x[3]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_x_reg[3]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_3_ ( .D(
        Inst_Gf16_mul2_Canright2_x[4]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_x_reg[4]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_4_ ( .D(
        Inst_Gf16_mul2_Canright2_y[1]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_y_reg[1]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_5_ ( .D(
        Inst_Gf16_mul2_Canright2_y[2]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_y_reg[2]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_6_ ( .D(
        Inst_Gf16_mul2_Canright2_y[3]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_y_reg[3]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_7_ ( .D(
        Inst_Gf16_mul2_Canright2_y[4]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_y_reg[4]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_8_ ( .D(
        Inst_Gf16_mul2_Canright2_z[1]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_z_reg[1]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_9_ ( .D(
        Inst_Gf16_mul2_Canright2_z[2]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_z_reg[2]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_10_ ( .D(
        Inst_Gf16_mul2_Canright2_z[3]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_z_reg[3]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_11_ ( .D(
        Inst_Gf16_mul2_Canright2_z[4]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_z_reg[4]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_12_ ( .D(
        Inst_Gf16_mul2_Canright2_t[1]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_t_reg[1]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_13_ ( .D(
        Inst_Gf16_mul2_Canright2_t[2]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_t_reg[2]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_14_ ( .D(
        Inst_Gf16_mul2_Canright2_t[3]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_t_reg[3]), .QN() );
  DFF_X1 Inst_Gf16_mul2_Canright2_GEN_reg_s_current_state_reg_15_ ( .D(
        Inst_Gf16_mul2_Canright2_t[4]), .CK(clk), .Q(
        Inst_Gf16_mul2_Canright2_t_reg[4]), .QN() );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst0_U1 ( 
        .A(Inst_Gf16_mul2_Canright2_x_reg[1]), .B(
        Inst_Gf16_mul2_Canright2_x_reg[2]), .Z(dcba1_out[0]) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst1_U1 ( 
        .A(Inst_Gf16_mul2_Canright2_x_reg[3]), .B(
        Inst_Gf16_mul2_Canright2_x_reg[4]), .Z(dcba2_out[0]) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst2_U1 ( 
        .A(Inst_Gf16_mul2_Canright2_y_reg[1]), .B(
        Inst_Gf16_mul2_Canright2_y_reg[2]), .Z(dcba1_out[1]) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst3_U1 ( 
        .A(Inst_Gf16_mul2_Canright2_y_reg[3]), .B(
        Inst_Gf16_mul2_Canright2_y_reg[4]), .Z(dcba2_out[1]) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst4_U1 ( 
        .A(Inst_Gf16_mul2_Canright2_z_reg[1]), .B(
        Inst_Gf16_mul2_Canright2_z_reg[2]), .Z(dcba1_out[2]) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst5_U1 ( 
        .A(Inst_Gf16_mul2_Canright2_z_reg[3]), .B(
        Inst_Gf16_mul2_Canright2_z_reg[4]), .Z(dcba2_out[2]) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst6_U1 ( 
        .A(Inst_Gf16_mul2_Canright2_t_reg[1]), .B(
        Inst_Gf16_mul2_Canright2_t_reg[2]), .Z(dcba1_out[3]) );
  XOR2_X1 Inst_Gf16_mul2_Canright2_Inst_Gf6_sq_scl_mul_Canright_L_XORInst7_U1 ( 
        .A(Inst_Gf16_mul2_Canright2_t_reg[3]), .B(
        Inst_Gf16_mul2_Canright2_t_reg[4]), .Z(dcba2_out[3]) );
endmodule

